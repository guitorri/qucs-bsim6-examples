* Modelcards from the BSIM6.1.0 benchmarks
* - This file contains the NMOS and PMOS modelcards
* - LEVEL and VERSION assigned to match Qucs current implementation
* - PMOS card was sed to UPPERCASE, qucsconv cannot map the paramter names otherwise
*

.model nmos NMOS LEVEL=6 VERSION=1.0
+LLONG =2E-06
+WWIDE =1E-05
+TYPE =1
+GEOMOD =0
+RGEOMOD =0
+COVMOD =1
+RDSMOD =0
+XL =-1.7E-08
+XW =1.1E-08
+LINT =0
+WINT =0
+DLC =0
+DWC =0
+TOXE =1.74E-09
+TOXP =1.7E-09
+NDEP =4.6E+23
+NSD =1E+26
+NGATE =8.5E+25
+VFB =-1.02
+EPSROX =3.9
+EPSRSUB =11.9
+NI0SUB =1.1E+16
+XJ =1.5E-07
+DMCG =0
+DMDG =0
+DMCGT =0
+CIT =1E-08
+CDSCD =0.001
+CDSCB =0
+CDSCBL =0.007
+CDSCBLEXP =1
+NFACTOR =0.002
+NFACTORL =2.1E-08
+NFACTORLEXP =6.264
+NDEPL1 =0.096
+NDEPLEXP1 =1
+NDEPL2 =-0.0032
+NDEPLEXP2 =2.05
+DVTP0 =7.5E-07
+DVTP1 =-4.4E-07
+NDEPW =-0.1548
+NDEPWEXP =0.7441
+NDEPWL =0
+NDEPWLEXP =0.2
+K2W =0
+GIDLMOD =1
+AGIDL =3.728E-08
+AGIDLL =-0.04815
+AGIDLW =-0.0341
+BGIDL =8.123E+09
+CGIDL =1.21E-06
+EGIDL =-2.952
+PHIN =0.05
+K2L =0.001636
+K2 =-0.014
+ETA0 =8.416E-06
+ETAB =-5.561E-05
+ETABEXP =2.155
+DSUB =3
+VSAT =6.4E+04
+VSATW =0.05
+VSATWEXP =1
+DELTA =0.15
+DELTAL =0.1
+DELTALEXP =1E-05
+U0 =0.04546
+ETAMOB =1.5
+U0L =0.025
+U0LEXP =0.95
+UA =0.4007
+UAW =0.05
+UAWEXP =1
+UAL =0.00475
+UALEXP =1.118
+EUW =-0.02
+EUWEXP =1
+EUL =0.001
+EULEXP =1
+EU =1.9
+UDL =1E-15
+UDLEXP =1
+UD =1.042E-05
+UCS =2
+UCW =0
+UCWEXP =1
+UC =1E-07
+UCL =2.5E+04
+UCLEXP =1
+PCLM =0.15
+PCLML =0.01
+PCLMLEXP =0.4
+PCLMG =0
+PSCBE1 =5
+PSCBE2 =1.29E-12
+PDITS =0
+PDITSL =0
+PDITSD =0
+RSWMIN =0
+RSW =100
+RDWMIN =0
+RDW =100
+RDSW =20
+RDSWMIN =0
+PRWG =1
+PRWB =0
+WR =1
+RSH =0
+PDIBLCB =0
+PDIBLC =0.01
+PDIBLCL =1E-05
+PDIBLCLEXP =1E-06
+PVAG =0
+PTWG =0.2
+PTWGL =3E+04
+PTWGLEXP =5E-06
+FPROUT =0
+CF =0
+CFRCOEFF =1
+CGSO =2.5E-10
+CGDO =2.5E-10
+CGSL =1.2E-10
+CGDL =1.2E-10
+CKAPPAS =1.25
+CKAPPAD =1.25
+CGBO =0
+ADOS =0
+BDOS =1
+QM0 =0.001
+ETAQM =0.54
+NDEPCV =8E+23
+VFBCV =-0.95
+VSATCV =1E+05
+PCLMCV =0
+PSAT =0.46
+PSATL =6
+PSATLEXP =0.06
+TNFACTOR =0
+TETA0 =0
+UTE =-1.4
+UTEL =-0.001
+UA1 =-0.0011
+UA1L =0
+UC1 =0
+UD1 =0
+UD1L =0
+UCSTE =-0.005
+PRT =0
+AT =-0.05
+ATL =-0.1
+TDELTA =-0.0048
+PTWGT =-0.002
+PTWGTL =0.01
+KT1 =-0.115
+KT1EXP =1
+KT1L =1.286E-09
+KT2 =-0.003157
+K2LEXP =1.698
+K2WEXP =0.005
+TBGASUB =0
+IGCMOD =0
+IGBMOD =0
+AIGS=0.0136
+BIGS=0.00171
+CIGS=0.075
+AIGSL=0
+AIGD=0.0136
+BIGD=0.00171
+CIGD=0.075
+AIGDL=0
+AIGC=0.01285
+LAIGC=2.132E-06
+BIGC=0.0013
+CIGC=0.013
+AIGCL=-0.01227
+PIGCD=1
+PIGCDL=6.196
+AIGBINV=0.015
+BIGBINV=0.000949
+CIGBINV=0.006
+EIGBINV=1.1
+NIGBINV=3
+AIGBACC=0.01751
+BIGBACC=8.307
+CIGBACC=-898.7
+NIGBACC=1
+LPSAT=0
+WPSAT=0
+PPSAT=0
+PSATB=0
+PSATX=3
+WVSAT=0
+PVSAT=0
+WPTWG=0
+PPTWG=0
+TNOM=25
+WDVTP0=0
+WDVTP1=0
+LUTE=0.04574
+LUA1=8.365E-05
+LAT=0
+DVTP2=0
+DVTP3=0
+DVTP4=0
+DVTP5=0
+VSATL=1350
+VSATLEXP=0.00033


.model pmos PMOS LEVEL=6 VERSION=1.0
+TOXE    = 2.34E-009
+TOXP    = 1.925E-009
+DTOX    = 0
+EPSROX  = 3.9
+TNOM    = 25
+XL      = 0
+XW      = 0
+LINT    = 0
+LLONG   = 1000000
+LL      = 0
+LW      = 0
+LWL     = 0
+LLN     = 1
+LWN     = 1
+WINT    = -9.0134104E-009
+WL      = 0
+WW      = 0
+WWL     = 0
+WLN     = 1
+WWN     = 1
+WWIDE   = 1000000
+DLC     = 0
+LLC     = 0
+LWC     = 0
+LWLC    = 0
+DWC     = 0
+WLC     = 0
+WWC     = 0
+WWLC    = 0
+GEOMOD  = 0
+RGEOMOD = 0
+RGATEMOD= 0
+RBODYMOD= 0
+IGCMOD  = 0
+IGBMOD  = 0
+COVMOD  = 1
+RDSMOD  = 0
+GIDLMOD = 0
+TNOIMOD = 0
+GMIN    = 1E-012
+JSS     = 0.0001
+JSD     = 0.0001
+JSWS    = 0
+JSWD    = 0
+JSWGS   = 0
+JSWGD   = 0
+NJS     = 1
+NJD     = 1
+IJTHSFWD= 0.1
+IJTHDFWD= 0.1
+IJTHSREV= 0.1
+IJTHDREV= 0.1
+BVS     = 10
+BVD     = 10
+XJBVS   = 1
+XJBVD   = 1
+JTSS    = 0
+JTSD    = 0
+JTSSWS  = 0
+JTSSWD  = 0
+JTSSWGS = 0
+JTSSWGD = 0
+JTWEFF  = 0
+NJTS    = 20
+NJTSD   = 20
+NJTSSW  = 20
+NJTSSWD = 20
+NJTSSWG = 20
+NJTSSWGD= 20
+VTSS    = 10
+VTSD    = 10
+VTSSWS  = 10
+VTSSWD  = 10
+VTSSWGS = 10
+VTSSWGD = 10
+CJS     = 0.0005
+CJD     = 0.0005
+CJSWS   = 5E-010
+CJSWD   = 5E-010
+CJSWGS  = 0
+CJSWGD  = 0
+PBS     = 1
+PBD     = 1
+PBSWS   = 1
+PBSWD   = 1
+PBSWGS  = 1
+PBSWGD  = 1
+MJS     = 0.5
+MJD     = 0.5
+MJSWS   = 0.33
+MJSWD   = 0.33
+MJSWGS  = 0.33
+MJSWGD  = 0.33
+TPB     = 0
+TCJ     = 0
+TPBSW   = 0
+TCJSW   = 0
+TPBSWG  = 0
+TCJSWG  = 0
+XTIS    = 3
+XTID    = 3
+XTSS    = 0.02
+XTSD    = 0.02
+XTSSWS  = 0.02
+XTSSWD  = 0.02
+XTSSWGS = 0.02
+XTSSWGD = 0.02
+TNJTS   = 0
+TNJTSD  = 0
+TNJTSSW = 0
+TNJTSSWD= 0
+TNJTSSWG= 0
+TNJTSSWGD= 0
+NOIA    = 6.25E+040
+NOIB    = 3.125E+025
+NOIC    = 8.75E+008
+EM      = 41000000
+EF      = 1
+LINTNOI = 0
+NTNOI   = 1
+TNOIA   = 0
+TNOIB   = 0
+TNOIC   = 0
+RNOIA   = 0.577
+RNOIB   = 0.5164
+RNOIC   = 0.395
+DWJ     = 0
+DMCG    = 0
+DMCI    = 0
+DMDG    = 0
+DMCGT   = 0
+XGW     = 0
+XGL     = 0
+GBMIN   = 1E-012
+RSHG    = 0.1
+RBPB    = 50
+RBPD    = 50
+RBPS    = 50
+RBDB    = 50
+RBSB    = 50
+RBPS0   = 50
+RBPSL   = 0
+RBPSW   = 0
+RBPSNF  = 0
+RBPD0   = 50
+RBPDL   = 0
+RBPDW   = 0
+RBPDNF  = 0
+RBPBX0  = 100
+RBPBXL  = 0
+RBPBXW  = 0
+RBPBXNF = 0
+RBPBY0  = 100
+RBPBYL  = 0
+RBPBYW  = 0
+RBPBYNF = 0
+RBSBX0  = 100
+RBSBY0  = 100
+RBDBX0  = 100
+RBDBY0  = 100
+RBSDBXL = 0
+RBSDBXW = 0
+RBSDBXNF= 0
+RBSDBYL = 0
+RBSDBYW = 0
+RBSDBYNF= 0
+XRCRG1  = 12
+XRCRG2  = 1
+NGCON   = 1
+NDEP    = 8.062E+023
+NDEPL1  = 1.2139
+NDEPLEXP1= 1.9088
+NDEPL2  = -1.1825
+NDEPLEXP2= 1.9173
+NDEPW   = 0.065035
+NDEPWEXP= 0.48882
+NDEPWL  = 0.00040893
+NDEPWLEXP= 1.3273
+EASUB   = 4.05
+NI0SUB  = 1.1E+016
+BG0SUB  = 1.17
+EPSRSUB = 11.9
+XJ      = 1.5E-007
+VFB     = -1.2108
+VFBSDOFF= 0
+NSD     = 1E+026
+DVTP0   = 1.8335E-007
+DVTP1   = 220.59
+DVTP2   = 9.6351E-010
+DVTP3   = 0.89017
+DVTP4   = 98.728
+DVTP5   = 5.1435E-017
+PHIN    = 0.045
+ETA0    = 0.0051075
+ETAB    = -0.010908157
+ETABEXP = 0.09999
+DSUB    = 1.0667
+K2      = -0.093146
+K2L     = 0.065574
+K2LEXP  = 0.79778
+K2W     = 0.030809
+K2WEXP  = 0.87253
+CIT     = 1.0136148E-005
+CDSCD   = 0.0011509049
+CDSCDL  = -0.00048388809
+CDSCDLEXP= 0.13963388
+CDSCB   = 9.9995516E-006
+CDSCBL  = 1.4756534E-009
+CDSCBLEXP= 1
+NFACTOR = 0.0017201
+NFACTORL= 1.7832E-006
+NFACTORLEXP= 0.99988
+NFACTORW= 0.11149
+NFACTORWEXP= 0.8993
+NFACTORWL= -0.01386
+U0      = 0.04004
+U0L     = 0.58676
+U0LEXP  = 0.11151
+ETAMOB  = 4.0947
+UA      = 0.4298
+UAL     = -0.0087246
+UALEXP  = 1.3647
+UAW     = 0.11575
+UAWEXP  = 0.4385
+UAWL    = -7.027E-005
+EU      = 1.3371
+EUL     = 0.0021948
+EULEXP  = 1.4769
+EUW     = -0.0031666
+EUWEXP  = 1.9366
+EUWL    = -0.00013929
+UD      = 0.0093995
+UDL     = 0.067484
+UDLEXP  = 0.099452
+UCS     = 0.9999
+UC      = 4.91E-006
+UCL     = 0.001096
+UCLEXP  = 0.0015937
+VSAT    = 9609100
+VSATL   = 6.8282
+VSATLEXP= 0.086396
+VSATW   = 0.016834
+VSATWEXP= 3.0172
+VSATCVL = 0
+VSATCVLEXP= 1
+VSATCVW = 0
+VSATCVWEXP= 1
+DELTA   = 0.1779
+DELTAL  = 0.1269
+DELTALEXP= 0.18156
+PCLM    = 0
+PCLML   = 0
+PCLMLEXP= 1E-013
+PCLMG   = 0
+PCLMCVL = 0
+PCLMCVLEXP= 1
+PSCBE1  = 4.24E+008
+PSCBE2  = 1E-008
+PDITS   = 0.85536
+PDITSL  = 8473.9
+PDITSD  = 0
+PDIBLC  = 0.005
+PDIBLCL = 0
+PDIBLCLEXP= 1
+PDIBLCB = -0.49995
+PVAG    = 1
+FPROUT  = 0
+FPROUTL = 0
+FPROUTLEXP= 1
+PTWG    = 0.09999
+PTWGL   = 0.069993
+PTWGLEXP= 0.0009999
+PSAT    = 1E-013
+PSATL   = 0
+PSATLEXP= 1
+PSATB   = 0.9999
+PSATX   = 1E-013
+RSH     = 0
+PRWG    = 1
+PRWB    = 0.010098993
+PRWBL   = 0.00070000265
+PRWBLEXP= 1
+WR      = 1
+RSWMIN  = 0
+RSW     = 10
+RSWL    = 0
+RSWLEXP = 1
+RDWMIN  = 0
+RDW     = 10
+RDWL    = 0
+RDWLEXP = 1
+RDSWMIN = 0
+RDSW    = 0
+RDSWL   = 0.0007
+RDSWLEXP= 1E-007
+ALPHA0  = 0
+ALPHA0L = 0
+ALPHA0LEXP= 1
+BETA0   = 0
+AGIDL   = 0
+AGIDLL  = 0
+AGIDLW  = 0
+BGIDL   = 2.3E+009
+CGIDL   = 0.5
+EGIDL   = 0.8
+AGISL   = 0
+AGISLL  = 0
+AGISLW  = 0
+BGISL   = 2.3E+009
+CGISL   = 0.5
+EGISL   = 0.00171
+AIGBACC = 0.00171
+BIGBACC = 0.00171
+CIGBACC = 0.075
+NIGBACC = 1
+AIGBINV = 0.0111
+BIGBINV = 0.000949
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC    = 0.0136
+AIGCL   = 3
+AIGCW   = 0.0136
+BIGC    = 0.00171
+CIGC    = 0.075
+AIGS    = 0.0136
+AIGSL   = 0.075
+AIGSW   = 0.0136
+AIGD    = 0.0136
+AIGDL   = 0
+AIGDW   = 0.0136
+BIGS    = 0.00171
+BIGD    = 0.00171
+CIGS    = 0.075
+CIGD    = 0.075
+TOXREF  = 0.075
+NTOX    = 1
+POXEDGE = 1
+PIGCD   = 1
+PIGCDL  = 1
+NDEPCV = 4.598E+23
+NDEPCVL1= 0
+NDEPCVLEXP1= 1
+NDEPCVL2= 0
+NDEPCVLEXP2= 2
+NDEPCVW = 0
+NDEPCVWEXP= 1
+NDEPCVWL= 0
+NDEPCVWLEXP= 1
+NGATE   = 7.764E+25
+CF      = 0
+CFRCOEFF= 1
+CGSO    = 187.0E-12
+CGDO    = 187.0E-12
+CGBO    = 0
+CGSL    = 130.0E-12
+CGDL    = 130.0E-12
+CKAPPAS = 1.6
+CKAPPAD = 1.6
+ADOS    = 221.4
+BDOS    = 1.350
+QM0     = 405.7E-6
+ETAQM   = 848.5E-3
+VFBCV   = -996.0E-3
+VFBCVL  = 0
+VFBCVLEXP= 1
+VFBCVW  = 0
+VFBCVWEXP= 1
+VFBCVWL = 0
+VFBCVWLEXP= 1
+TBGASUB = 0.000473
+TBGBSUB = 636
+TDELTA  = 0
+PTWGT   = 0
+IIT     = 0
+TGIDL   = 0
+IGT     = 0
+KT1     = -0.11
+KT1L    = 0
+KT2     = 0.022
+KT1EXP  = 1
+UTE     = -1.5
+UA1     = 0.001
+UD1     = 0
+UC1     = -5.6E-011
+UCSTE   = -0.004775
+PRT     = 0
+AT      = -0.00156
+SCA     = 0
+SCB     = 0
+SCC     = 0
+SC      = 0
+KU0WE   = 0
+KVTH0WE = 0
+K2WE    = 0
+WEB     = 0
+WEC     = 0
+SCREF   = 1E-006
+SA      = 0
+SB      = 0
+SD      = 0
+SAREF   = 1E-006
+SBREF   = 1E-006
+WLOD    = 0
+KVSAT   = 0
+KU0     = 0
+TKU0    = 0
+LKU0    = 0
+WKU0    = 0
+PKU0    = 0
+LLODKU0 = 0
+WLODKU0 = 0
+KVTH0   = 0
+LKVTH0  = 0
+WKVTH0  = 0
+PKVTH0  = 0
+LLODVTH = 0
+WLODVTH = 0
+STK2    = 0
+LODK2   = 1
+STETA0  = 0
+LODETA0 = 1


.END

